package test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import simple_env_pkg::simple_env;
    import simple_agent_pkg::*;

    `include "base_test.sv"
    `include "simple_test.sv"

endpackage
