package simple_env_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import simple_agent_pkg::*;

    `include "simple_env.sv"
endpackage : simple_env_pkg