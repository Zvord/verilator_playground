package test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import simple_env_pkg::simple_env;

    `include "base_test.sv"

endpackage