class item extends uvm_sequence_item;
endclass