package simple_agent_pkg;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "simple_item.sv"
    `include "simple_sequencer.sv"
    `include "simple_driver.sv"
    `include "simple_monitor.sv"
    `include "simple_agent.sv"
    `include "simple_sequence.sv"
endpackage